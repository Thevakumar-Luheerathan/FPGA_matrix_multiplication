module control_unit_test();

	control_unit cu1();

endmodule